:insert

/*
*******************************************************************************
* File:        upsAgsIgrReplayCheckDtlsEpochTest.sv
*
* Author:       Shekhar Agrawal <sheagraw@cisco.com>
* Created:      Mar 17, 2010
* Language:     SystemVerilog
*
* Copyright 2009 Cisco Systems, Inc., All Rights Reserved.
* Cisco Systems Confidential
*
*******************************************************************************
* Description:
********************************************************************************
*/


.
